library ieee;
use ieee.std_logic_1164.all;

package types is
--  subtype row_range is natural range 0 to 7;
--  subtype col_range is natural range 7 downto 0;

end package;
